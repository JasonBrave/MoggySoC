module cpu_subsys_sram (
    input logic			clk,
    input logic			rst_n,
    input logic			mem_valid,
    input logic [29:0]	mem_addr,
	input logic			mem_write,
    input logic [31:0]	mem_wdata,
    input logic [3:0]	mem_wstrb,
    output logic [31:0]	mem_rdata,
    output logic		mem_ready);

    logic [31:0] mem [16384-1:0];

    always_ff @(posedge clk) begin
        if(mem_valid) begin
			if(mem_write) begin
				if(mem_wstrb[0]) mem[mem_addr[15:2]][7:0] <= mem_wdata[7:0];
				if(mem_wstrb[1]) mem[mem_addr[15:2]][15:8] <= mem_wdata[15:8];
				if(mem_wstrb[2]) mem[mem_addr[15:2]][23:16] <= mem_wdata[23:16];
				if(mem_wstrb[3]) mem[mem_addr[15:2]][31:24] <= mem_wdata[31:24];
			end

			mem_rdata <= mem[mem_addr[15:2]];
			mem_ready <= 1'b1;
        end else begin
			mem_ready <= 1'b0;
		end
    end

endmodule // cpu_subsys_sram
