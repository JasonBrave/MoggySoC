module interconnect_subsys_tb;
endmodule
